library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package Common is
    type CHAR_ARRAY is array (integer range<>) of std_logic_vector(7 downto 0);
end Common;

package body Common is
   -- subprogram bodies here
end Common;